module main

struct User {
	id    int
	name string
	phone  string
}